*tristate

.SUBCKT TI IN ZN EN VDD VSS
*M_i Drain Gate Source Bulk
M_i_0 1 A VSS VSS NMOS W=0.415000U L=0.050000U
M_i_2 ZN EN 1 VSS NMOS W=0.415000U L=0.050000U

M_i_3 2 ENB ZN VDD PMOS W=0.630000U L=0.050000U
M_i_1 VDD A 2 VDD PMOS W=0.630000U L=0.050000U

M_i_4 A IN VDD VDD PMOS W=0.630000U L=0.050000U
M_i_5 A IN VSS VSS NMOS W=0.630000U L=0.050000U

M_i_6 ENB EN VDD VDD PMOS W=0.630000U L=0.050000U
M_i_7 ENB EN VSS VSS NMOS W=0.630000U L=0.050000U
.ENDS 
