.include '45nm_LP.pm'

.SUBCKT PT A Y EN ENB
*M_i Drain Gate Source Bulk
M_i_0 Y EN A A NMOS W=0.415000U L=0.050000U
M_i_2 Y ENB A A PMOS W=0.415000U L=0.050000U
.ENDS 

