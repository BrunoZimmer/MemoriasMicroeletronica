*Tristate inverter

.SUBCKT TI A ZN EN ENB VDD VSS 
*M_i Drain Gate Source Bulk
M_i_0 1 A VSS VSS NMOS W=0.415000U L=0.050000U
M_i_2 ZN EN 1 VSS NMOS W=0.415000U L=0.050000U

M_i_3 2 ENB ZN VDD PMOS W=0.630000U L=0.050000U
M_i_1 VDD A 2 VDD PMOS W=0.630000U L=0.050000U
.ENDS 

